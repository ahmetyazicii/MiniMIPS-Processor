module and32(
	input [31:0]A,
	input [31:0]B,
	output [31:0]R
	);

	
	// and 32 bits one by one
	and and31(R[31],A[31],B[31]);
	and and30(R[30],A[30],B[30]);
	and and29(R[29],A[29],B[29]);
	and and28(R[28],A[28],B[28]);
	and and27(R[27],A[27],B[27]);
	and and26(R[26],A[26],B[26]);
	and and25(R[25],A[25],B[25]);
	and and24(R[24],A[24],B[24]);
	and and23(R[23],A[23],B[23]);
	and and22(R[22],A[22],B[22]);
	and and21(R[21],A[21],B[21]);
	and and20(R[20],A[20],B[20]);
	and and19(R[19],A[19],B[19]);
	and and18(R[18],A[18],B[18]);
	and and17(R[17],A[17],B[17]);
	and and16(R[16],A[16],B[16]);
	and and15(R[15],A[15],B[15]);
	and and14(R[14],A[14],B[14]);
	and and13(R[13],A[13],B[13]);
	and and12(R[12],A[12],B[12]);
	and and11(R[11],A[11],B[11]);
	and and10(R[10],A[10],B[10]);
	and and9(R[9],A[9],B[9]);
	and and8(R[8],A[8],B[8]);
	and and7(R[7],A[7],B[7]);
	and and6(R[6],A[6],B[6]);
	and and5(R[5],A[5],B[5]);
	and and4(R[4],A[4],B[4]);
	and and3(R[3],A[3],B[3]);
	and and2(R[2],A[2],B[2]);
	and and1(R[1],A[1],B[1]);
	and and0(R[0],A[0],B[0]);
	

endmodule