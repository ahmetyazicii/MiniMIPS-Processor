module or32(
	input [31:0]A,
	input [31:0]B,
	output [31:0]R
	);

	// or 32 bits one by one
	or or31(R[31],A[31],B[31]);
	or or30(R[30],A[30],B[30]);
	or or29(R[29],A[29],B[29]);
	or or28(R[28],A[28],B[28]);
	or or27(R[27],A[27],B[27]);
	or or26(R[26],A[26],B[26]);
	or or25(R[25],A[25],B[25]);
	or or24(R[24],A[24],B[24]);
	or or23(R[23],A[23],B[23]);
	or or22(R[22],A[22],B[22]);
	or or21(R[21],A[21],B[21]);
	or or20(R[20],A[20],B[20]);
	or or19(R[19],A[19],B[19]);
	or or18(R[18],A[18],B[18]);
	or or17(R[17],A[17],B[17]);
	or or16(R[16],A[16],B[16]);
	or or15(R[15],A[15],B[15]);
	or or14(R[14],A[14],B[14]);
	or or13(R[13],A[13],B[13]);
	or or12(R[12],A[12],B[12]);
	or or11(R[11],A[11],B[11]);
	or or10(R[10],A[10],B[10]);
	or or9(R[9],A[9],B[9]);
	or or8(R[8],A[8],B[8]);
	or or7(R[7],A[7],B[7]);
	or or6(R[6],A[6],B[6]);
	or or5(R[5],A[5],B[5]);
	or or4(R[4],A[4],B[4]);
	or or3(R[3],A[3],B[3]);
	or or2(R[2],A[2],B[2]);
	or or1(R[1],A[1],B[1]);
	or or0(R[0],A[0],B[0]);
	

endmodule