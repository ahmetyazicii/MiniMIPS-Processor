module nor32(
	input [31:0]A,
	input [31:0]B,
	output [31:0]R
	);

	// nor 32 bits one by one
	nor nor31(R[31],A[31],B[31]);
	nor nor30(R[30],A[30],B[30]);
	nor nor29(R[29],A[29],B[29]);
	nor nor28(R[28],A[28],B[28]);
	nor nor27(R[27],A[27],B[27]);
	nor nor26(R[26],A[26],B[26]);
	nor nor25(R[25],A[25],B[25]);
	nor nor24(R[24],A[24],B[24]);
	nor nor23(R[23],A[23],B[23]);
	nor nor22(R[22],A[22],B[22]);
	nor nor21(R[21],A[21],B[21]);
	nor nor20(R[20],A[20],B[20]);
	nor nor19(R[19],A[19],B[19]);
	nor nor18(R[18],A[18],B[18]);
	nor nor17(R[17],A[17],B[17]);
	nor nor16(R[16],A[16],B[16]);
	nor nor15(R[15],A[15],B[15]);
	nor nor14(R[14],A[14],B[14]);
	nor nor13(R[13],A[13],B[13]);
	nor nor12(R[12],A[12],B[12]);
	nor nor11(R[11],A[11],B[11]);
	nor nor10(R[10],A[10],B[10]);
	nor nor9(R[9],A[9],B[9]);
	nor nor8(R[8],A[8],B[8]);
	nor nor7(R[7],A[7],B[7]);
	nor nor6(R[6],A[6],B[6]);
	nor nor5(R[5],A[5],B[5]);
	nor nor4(R[4],A[4],B[4]);
	nor nor3(R[3],A[3],B[3]);
	nor nor2(R[2],A[2],B[2]);
	nor nor1(R[1],A[1],B[1]);
	nor nor0(R[0],A[0],B[0]);
	

endmodule